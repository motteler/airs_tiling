netcdf airs_tiling {
dimensions:
	obs = 12150 ;
	wnum = 2645 ;
variables:
	double tai93(obs) ;
		tai93:valid_range = -2934835217., 3376598410. ;
		string tai93:long_name = "earth view FOV midtime" ;
		tai93:_FillValue = 9.96920996838687e+36 ;
		string tai93:coverage_content_type = "referenceInformation" ;
		string tai93:standard_name = "time" ;
		string tai93:units = "seconds since 1993-01-01 00:00" ;
		string tai93:description = "earth view observation midtime for each FOV" ;
		string tai93:AIRS_HDF_name = "Time" ;
	float lat(obs) ;
		lat:valid_range = -90.f, 90.f ;
		string lat:long_name = "latitude" ;
		lat:_FillValue = 9.96921e+36f ;
		string lat:bounds = "lat_bnds" ;
		string lat:coverage_content_type = "referenceInformation" ;
		string lat:standard_name = "latitude" ;
		string lat:units = "degrees_north" ;
		string lat:description = "latitude of FOV center" ;
		string lat:AIRS_HDF_name = "Latitude" ;
	float lon(obs) ;
		lon:valid_range = -180.f, 180.f ;
		string lon:long_name = "FOV longitude" ;
		lon:_FillValue = 9.96921e+36f ;
		string lon:bounds = "lon_bnds" ;
		string lon:coverage_content_type = "referenceInformation" ;
		string lon:standard_name = "longitude" ;
		string lon:units = "degrees_east" ;
		string lon:description = "longitude of FOV center" ;
		string lon:AIRS_HDF_name = "Longitude" ;
	float land_frac(obs) ;
		land_frac:valid_range = 0.f, 1.f ;
		string land_frac:long_name = "land fraction" ;
		string land_frac:coordinates = "lon lat" ;
		land_frac:_FillValue = 9.96921e+36f ;
		string land_frac:coverage_content_type = "referenceInformation" ;
		string land_frac:standard_name = "land_area_fraction" ;
		string land_frac:units = "1" ;
		string land_frac:description = "land fraction over the FOV" ;
		string land_frac:AIRS_HDF_name = "landFrac" ;
		string land_frac:cell_methods = "area: mean (beam-weighted)" ;
	float sol_zen(obs) ;
		sol_zen:valid_range = 0.f, 180.f ;
		string sol_zen:long_name = "solar zenith angle" ;
		string sol_zen:coordinates = "lon lat" ;
		sol_zen:_FillValue = 9.96921e+36f ;
		string sol_zen:coverage_content_type = "referenceInformation" ;
		string sol_zen:standard_name = "solar_zenith_angle" ;
		string sol_zen:units = "degree" ;
		string sol_zen:description = "solar zenith angle at the center of the FOV" ;
		string sol_zen:AIRS_HDF_name = "solzen" ;
	float sat_zen(obs) ;
		sat_zen:valid_range = 0.f, 180.f ;
		string sat_zen:long_name = "satellite zenith angle" ;
		string sat_zen:coordinates = "lon lat" ;
		sat_zen:_FillValue = 9.96921e+36f ;
		string sat_zen:coverage_content_type = "referenceInformation" ;
		string sat_zen:standard_name = "sensor_zenith_angle" ;
		string sat_zen:units = "degree" ;
		string sat_zen:description = "satellite zenith angle at the center of the FOV" ;
		string sat_zen:AIRS_HDF_name = "satzen" ;
	ubyte asc_flag(obs) ;
		asc_flag:valid_range = 0UB, 1UB ;
		string asc_flag:long_name = "ascending orbit flag" ;
		string asc_flag:coordinates = "subsat_lon subsat_lat" ;
		asc_flag:_FillValue = 255UB ;
		asc_flag:flag_values = 0UB, 1UB ;
		string asc_flag:coverage_content_type = "referenceInformation" ;
		string asc_flag:description = "ascending orbit flag: 1 if ascending, 0 descending" ;
		string asc_flag:AIRS_HDF_name = "scan_node_type" ;
		string asc_flag:flag_meanings = "descending ascending" ;
	float rad(obs, wnum) ;
		string rad:units = "mW/(m2 sr cm-1)" ;
		string rad:ancillary_variables = "rad_qc synth_frac chan_qc" ;
		string rad:long_name = "spectral radiance" ;
		string rad:standard_name = "toa_outgoing_radiance_per_unit_wavenumber" ;
		string rad:coordinates = "lon lat" ;
		string rad:description = "spectral radiance" ;
		rad:_FillValue = 9.96921e+36f ;
		string rad:coverage_content_type = "physicalMeasurement" ;
	byte rad_qc(obs) ;
		rad_qc:valid_range = 0b, 2b ;
		string rad_qc:long_name = "rad QC" ;
		string rad_qc:standard_name = "toa_outgoing_radiance_per_unit_wavenumber status_flag" ;
		string rad_qc:coordinates = "lon lat" ;
		string rad_qc:description = "rad QC flag" ;
		rad_qc:_FillValue = -1b ;
		string rad_qc:coverage_content_type = "qualityInformation" ;
		string rad_qc:flag_meanings = "Best Good Do_Not_Use" ;
		rad_qc:flag_values = 0b, 1b, 2b ;
	float synth_frac(wnum) ;
		string synth_frac:units = "1" ;
		synth_frac:valid_range = 0.f, 1.f ;
		string synth_frac:long_name = "Fraction synthesized" ;
		string synth_frac:description = "File mean fraction of signal that is attributed to synthesized AIRS Level-1C values" ;
		synth_frac:_FillValue = 9.96921e+36f ;
		string synth_frac:coverage_content_type = "qualityInformation" ;
	byte chan_qc(wnum) ;
		chan_qc:valid_range = 0b, 2b ;
		string chan_qc:long_name = "Channel QC" ;
		string chan_qc:standard_name = "toa_outgoing_radiance_per_unit_wavenumber status_flag" ;
		string chan_qc:description = "Quality of each channel." ;
		chan_qc:_FillValue = -1b ;
		string chan_qc:coverage_content_type = "qualityInformation" ;
		string chan_qc:flag_meanings = "Best Good Do_Not_Use" ;
		chan_qc:flag_values = 0b, 1b, 2b ;
	float nedn(wnum) ;
		string nedn:units = "mW/(m2 sr cm-1)" ;
		string nedn:long_name = "noise equivalent differential radiance" ;
		string nedn:description = "noise equivalent differential radiance" ;
		nedn:_FillValue = 9.96921e+36f ;
		string nedn:coverage_content_type = "qualityInformation" ;
	double wnum(wnum) ;
		string wnum:units = "cm-1" ;
		wnum:valid_range = 640., 2700. ;
		string wnum:long_name = "wavenumber" ;
		string wnum:standard_name = "sensor_band_central_radiation_wavenumber" ;
		string wnum:description = "wavenumber" ;
		wnum:_FillValue = 9.96920996838687e+36 ;
		string wnum:coverage_content_type = "auxiliaryInformation" ;
}
